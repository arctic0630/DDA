//memoria de instrucciones
module memins(
    input [31:0] fPC,
    output reg [31:0] ins
    );
    
    always @(*)
    begin
        casex(fPC)
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0000: ins = 32'b000000_00001_00010_00100_00000_100000; //suma
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0010: ins = 32'b000000_00001_00010_00100_00000_100010; //resta
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0011: ins = 32'b000000_00001_00010_00100_00000_100100; //and &
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0100: ins = 32'b000000_00001_00010_00100_00000_100101; //or
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0101: ins = 32'b000000_00001_00010_00100_00000_100110; //Xor
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0110: ins = 32'b000000_00001_00010_00100_00000_011000; //multiplicación
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX0111: ins = 32'b000100_00001_00010_0010000000000000; //branch
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX1000: ins = 32'b001000_00001_00010_0010000000000000; //desplazamiento
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX1001: ins = 32'b100011_00001_00010_0010000000000000; //load
            32'bXXXXXXXXXXXXXXXXXXXXXXXXXXXX1010: ins = 32'b001100_00001_00010_0010000000000000;
        endcase   
   end
endmodule     
